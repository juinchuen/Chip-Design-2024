module InputSignalRouter #(
    parameter D_WIDTH = 64,
    parameter LOG_2_WIDTH = 6
) (
    input logic [15:0] input_sig_Re [((D_WIDTH) - 1):0],
    input logic [15:0] input_sig_Im [((D_WIDTH) - 1):0],
    output logic [15:0] output_sig_Re [((D_WIDTH) - 1):0],
    output logic [15:0] output_sig_Im [((D_WIDTH) - 1):0]
);
    // Correctly route the input signal

    logic [15:0] fft_Re [((D_WIDTH) - 1):0];
    logic [15:0] fft_Im [((D_WIDTH) - 1):0];
	assign fft_Re[0] = input_sig_Re[0];
	assign fft_Im[0] = input_sig_Im[0];
	assign fft_Re[1] = input_sig_Re[32];
	assign fft_Im[1] = input_sig_Im[32];
	assign fft_Re[2] = input_sig_Re[16];
	assign fft_Im[2] = input_sig_Im[16];
	assign fft_Re[3] = input_sig_Re[48];
	assign fft_Im[3] = input_sig_Im[48];
	assign fft_Re[4] = input_sig_Re[8];
	assign fft_Im[4] = input_sig_Im[8];
	assign fft_Re[5] = input_sig_Re[40];
	assign fft_Im[5] = input_sig_Im[40];
	assign fft_Re[6] = input_sig_Re[24];
	assign fft_Im[6] = input_sig_Im[24];
	assign fft_Re[7] = input_sig_Re[56];
	assign fft_Im[7] = input_sig_Im[56];
	assign fft_Re[8] = input_sig_Re[4];
	assign fft_Im[8] = input_sig_Im[4];
	assign fft_Re[9] = input_sig_Re[36];
	assign fft_Im[9] = input_sig_Im[36];
	assign fft_Re[10] = input_sig_Re[20];
	assign fft_Im[10] = input_sig_Im[20];
	assign fft_Re[11] = input_sig_Re[52];
	assign fft_Im[11] = input_sig_Im[52];
	assign fft_Re[12] = input_sig_Re[12];
	assign fft_Im[12] = input_sig_Im[12];
	assign fft_Re[13] = input_sig_Re[44];
	assign fft_Im[13] = input_sig_Im[44];
	assign fft_Re[14] = input_sig_Re[28];
	assign fft_Im[14] = input_sig_Im[28];
	assign fft_Re[15] = input_sig_Re[60];
	assign fft_Im[15] = input_sig_Im[60];
	assign fft_Re[16] = input_sig_Re[2];
	assign fft_Im[16] = input_sig_Im[2];
	assign fft_Re[17] = input_sig_Re[34];
	assign fft_Im[17] = input_sig_Im[34];
	assign fft_Re[18] = input_sig_Re[18];
	assign fft_Im[18] = input_sig_Im[18];
	assign fft_Re[19] = input_sig_Re[50];
	assign fft_Im[19] = input_sig_Im[50];
	assign fft_Re[20] = input_sig_Re[10];
	assign fft_Im[20] = input_sig_Im[10];
	assign fft_Re[21] = input_sig_Re[42];
	assign fft_Im[21] = input_sig_Im[42];
	assign fft_Re[22] = input_sig_Re[26];
	assign fft_Im[22] = input_sig_Im[26];
	assign fft_Re[23] = input_sig_Re[58];
	assign fft_Im[23] = input_sig_Im[58];
	assign fft_Re[24] = input_sig_Re[6];
	assign fft_Im[24] = input_sig_Im[6];
	assign fft_Re[25] = input_sig_Re[38];
	assign fft_Im[25] = input_sig_Im[38];
	assign fft_Re[26] = input_sig_Re[22];
	assign fft_Im[26] = input_sig_Im[22];
	assign fft_Re[27] = input_sig_Re[54];
	assign fft_Im[27] = input_sig_Im[54];
	assign fft_Re[28] = input_sig_Re[14];
	assign fft_Im[28] = input_sig_Im[14];
	assign fft_Re[29] = input_sig_Re[46];
	assign fft_Im[29] = input_sig_Im[46];
	assign fft_Re[30] = input_sig_Re[30];
	assign fft_Im[30] = input_sig_Im[30];
	assign fft_Re[31] = input_sig_Re[62];
	assign fft_Im[31] = input_sig_Im[62];
	assign fft_Re[32] = input_sig_Re[1];
	assign fft_Im[32] = input_sig_Im[1];
	assign fft_Re[33] = input_sig_Re[33];
	assign fft_Im[33] = input_sig_Im[33];
	assign fft_Re[34] = input_sig_Re[17];
	assign fft_Im[34] = input_sig_Im[17];
	assign fft_Re[35] = input_sig_Re[49];
	assign fft_Im[35] = input_sig_Im[49];
	assign fft_Re[36] = input_sig_Re[9];
	assign fft_Im[36] = input_sig_Im[9];
	assign fft_Re[37] = input_sig_Re[41];
	assign fft_Im[37] = input_sig_Im[41];
	assign fft_Re[38] = input_sig_Re[25];
	assign fft_Im[38] = input_sig_Im[25];
	assign fft_Re[39] = input_sig_Re[57];
	assign fft_Im[39] = input_sig_Im[57];
	assign fft_Re[40] = input_sig_Re[5];
	assign fft_Im[40] = input_sig_Im[5];
	assign fft_Re[41] = input_sig_Re[37];
	assign fft_Im[41] = input_sig_Im[37];
	assign fft_Re[42] = input_sig_Re[21];
	assign fft_Im[42] = input_sig_Im[21];
	assign fft_Re[43] = input_sig_Re[53];
	assign fft_Im[43] = input_sig_Im[53];
	assign fft_Re[44] = input_sig_Re[13];
	assign fft_Im[44] = input_sig_Im[13];
	assign fft_Re[45] = input_sig_Re[45];
	assign fft_Im[45] = input_sig_Im[45];
	assign fft_Re[46] = input_sig_Re[29];
	assign fft_Im[46] = input_sig_Im[29];
	assign fft_Re[47] = input_sig_Re[61];
	assign fft_Im[47] = input_sig_Im[61];
	assign fft_Re[48] = input_sig_Re[3];
	assign fft_Im[48] = input_sig_Im[3];
	assign fft_Re[49] = input_sig_Re[35];
	assign fft_Im[49] = input_sig_Im[35];
	assign fft_Re[50] = input_sig_Re[19];
	assign fft_Im[50] = input_sig_Im[19];
	assign fft_Re[51] = input_sig_Re[51];
	assign fft_Im[51] = input_sig_Im[51];
	assign fft_Re[52] = input_sig_Re[11];
	assign fft_Im[52] = input_sig_Im[11];
	assign fft_Re[53] = input_sig_Re[43];
	assign fft_Im[53] = input_sig_Im[43];
	assign fft_Re[54] = input_sig_Re[27];
	assign fft_Im[54] = input_sig_Im[27];
	assign fft_Re[55] = input_sig_Re[59];
	assign fft_Im[55] = input_sig_Im[59];
	assign fft_Re[56] = input_sig_Re[7];
	assign fft_Im[56] = input_sig_Im[7];
	assign fft_Re[57] = input_sig_Re[39];
	assign fft_Im[57] = input_sig_Im[39];
	assign fft_Re[58] = input_sig_Re[23];
	assign fft_Im[58] = input_sig_Im[23];
	assign fft_Re[59] = input_sig_Re[55];
	assign fft_Im[59] = input_sig_Im[55];
	assign fft_Re[60] = input_sig_Re[15];
	assign fft_Im[60] = input_sig_Im[15];
	assign fft_Re[61] = input_sig_Re[47];
	assign fft_Im[61] = input_sig_Im[47];
	assign fft_Re[62] = input_sig_Re[31];
	assign fft_Im[62] = input_sig_Im[31];
	assign fft_Re[63] = input_sig_Re[63];
	assign fft_Im[63] = input_sig_Im[63];
	assign output_sig_Re = fft_Re;
	assign output_sig_Im = fft_Im;
endmodule
