`define ReW0 12'd2048
`define ReW1or63 12'd2040
`define ReW2or62 12'd2008
`define ReW3or61 12'd1960
`define ReW4or60 12'd1896
`define ReW5or59 12'd1808
`define ReW6or58 12'd1704
`define ReW7or57 12'd1584
`define ReW8or56 12'd1448
`define ReW9or55 12'd1296
`define ReW10or54 12'd1136
`define ReW11or53 12'd968
`define ReW12or52 12'd784
`define ReW13or51 12'd592
`define ReW14or50 12'd400
`define ReW15or49 12'd200
`define ReW16or48 12'd0
`define ReW17or47 12'd-200
`define ReW18or46 12'd-400
`define ReW19or45 12'd-592
`define ReW20or44 12'd-784
`define ReW21or43 12'd-968
`define ReW22or42 12'd-1136
`define ReW23or41 12'd-1296
`define ReW24or40 12'd-1448
`define ReW25or39 12'd-1584
`define ReW26or38 12'd-1704
`define ReW27or37 12'd-1808
`define ReW28or36 12'd-1896
`define ReW29or35 12'd-1960
`define ReW30or34 12'd-2008
`define ReW31or33 12'd-2040
`define ReW32 12'd-2048
`define ImW0or32 = 12'd0
`define ImW1or31 = 12'd200
`define ImW2or30 = 12'd400
`define ImW3or29 = 12'd592
`define ImW4or28 = 12'd784
`define ImW5or27 = 12'd968
`define ImW6or26 = 12'd1136
`define ImW7or25 = 12'd1296
`define ImW8or24 = 12'd1448
`define ImW9or23 = 12'd1584
`define ImW10or22 = 12'd1704
`define ImW11or21 = 12'd1808
`define ImW12or20 = 12'd1896
`define ImW13or19 = 12'd1960
`define ImW14or18 = 12'd2008
`define ImW15or17 = 12'd2040
`define ImW16 = 12'd2048
`define ImW33or63 = 12'd-200
`define ImW34or62 = 12'd-400
`define ImW35or61 = 12'd-592
`define ImW36or60 = 12'd-784
`define ImW37or59 = 12'd-968
`define ImW38or58 = 12'd-1136
`define ImW39or57 = 12'd-1296
`define ImW40or56 = 12'd-1448
`define ImW41or55 = 12'd-1584
`define ImW42or54 = 12'd-1704
`define ImW43or53 = 12'd-1808
`define ImW44or52 = 12'd-1896
`define ImW45or51 = 12'd-1960
`define ImW46or50 = 12'd-2008
`define ImW47or49 = 12'd-2040
`define ImW48 = 12'd-2048
