module InputSignalRouter #(
    parameter D_WIDTH = 64,
    parameter LOG_2_WIDTH = 6
) (
    input logic [1023:0] inputRe,
    input logic [1023:0] inputIm,
    output logic [1023:0] outputRe,
    output logic [1023:0] outputIm
);
    // Correctly route the input signal

    logic [1023:0] fftRe;
    logic [1023:0] fftIm;
	assign fftRe[0 +: 16] = inputRe[16 +: 15];
	assign fftIm[0 +: 16] = inputIm[16 +: 15];
	assign fftRe[1* 16 +: 16] = inputRe[32* 16 +: 16];
	assign fftIm[1* 16 +: 16] = inputIm[32* 16 +: 16];
	assign fftRe[2* 16 +: 16] = inputRe[16* 16 +: 16];
	assign fftIm[2* 16 +: 16] = inputIm[16* 16 +: 16];
	assign fftRe[3* 16 +: 16] = inputRe[48* 16 +: 16];
	assign fftIm[3* 16 +: 16] = inputIm[48* 16 +: 16];
	assign fftRe[4* 16 +: 16] = inputRe[8* 16 +:  16];
	assign fftIm[4* 16 +: 16] = inputIm[8* 16 +:  16];
	assign fftRe[5* 16 +: 16] = inputRe[40* 16 +: 16];
	assign fftIm[5* 16 +: 16] = inputIm[40* 16 +: 16];
	assign fftRe[6* 16 +: 16] = inputRe[24* 16 +: 16];
	assign fftIm[6* 16 +: 16] = inputIm[24* 16 +: 16];
	assign fftRe[7* 16 +: 16] = inputRe[56* 16 +: 16];
	assign fftIm[7* 16 +: 16] = inputIm[56* 16 +: 16];
	assign fftRe[8* 16 +: 16] = inputRe[4* 16 +: 16];
	assign fftIm[8* 16 +: 16] = inputIm[4* 16 +: 16];
	assign fftRe[9* 16 +: 16] = inputRe[36* 16 +: 16];
	assign fftIm[9* 16 +: 16] = inputIm[36* 16 +: 16];
	assign fftRe[10* 16 +: 16] = inputRe[20* 16 +: 16];
	assign fftIm[10* 16 +: 16] = inputIm[20* 16 +: 16];
	assign fftRe[11* 16 +: 16] = inputRe[52* 16 +: 16];
	assign fftIm[11* 16 +: 16] = inputIm[52* 16 +: 16];
	assign fftRe[12* 16 +: 16] = inputRe[12* 16 +: 16];
	assign fftIm[12* 16 +: 16] = inputIm[12* 16 +: 16];
	assign fftRe[13* 16 +: 16] = inputRe[44* 16 +: 16];
	assign fftIm[13* 16 +: 16] = inputIm[44* 16 +: 16];
	assign fftRe[14* 16 +: 16] = inputRe[28* 16 +: 16];
	assign fftIm[14* 16 +: 16] = inputIm[28* 16 +: 16];
	assign fftRe[15* 16 +: 16] = inputRe[60* 16 +: 16];
	assign fftIm[15* 16 +: 16] = inputIm[60* 16 +: 16];
	assign fftRe[16* 16 +: 16] = inputRe[2* 16 +: 16];
	assign fftIm[16* 16 +: 16] = inputIm[2* 16 +: 16];
	assign fftRe[17* 16 +: 16] = inputRe[34* 16 +: 16];
	assign fftIm[17* 16 +: 16] = inputIm[34* 16 +: 16];
	assign fftRe[18* 16 +: 16] = inputRe[18* 16 +: 16];
	assign fftIm[18* 16 +: 16] = inputIm[18* 16 +: 16];
	assign fftRe[19* 16 +: 16] = inputRe[50* 16 +: 16];
	assign fftIm[19* 16 +: 16] = inputIm[50* 16 +: 16];
	assign fftRe[20* 16 +: 16] = inputRe[10* 16 +: 16];
	assign fftIm[20* 16 +: 16] = inputIm[10* 16 +: 16];
	assign fftRe[21* 16 +: 16] = inputRe[42* 16 +: 16];
	assign fftIm[21* 16 +: 16] = inputIm[42* 16 +: 16];
	assign fftRe[22* 16 +: 16] = inputRe[26* 16 +: 16];
	assign fftIm[22* 16 +: 16] = inputIm[26* 16 +: 16];
	assign fftRe[23* 16 +: 16] = inputRe[58* 16 +: 16];
	assign fftIm[23* 16 +: 16] = inputIm[58* 16 +: 16];
	assign fftRe[24* 16 +: 16] = inputRe[6* 16 +: 16];
	assign fftIm[24* 16 +: 16] = inputIm[6* 16 +: 16];
	assign fftRe[25* 16 +: 16] = inputRe[38* 16 +: 16];
	assign fftIm[25* 16 +: 16] = inputIm[38* 16 +: 16];
	assign fftRe[26* 16 +: 16] = inputRe[22* 16 +: 16];
	assign fftIm[26* 16 +: 16] = inputIm[22* 16 +: 16];
	assign fftRe[27* 16 +: 16] = inputRe[54* 16 +: 16];
	assign fftIm[27* 16 +: 16] = inputIm[54* 16 +: 16];
	assign fftRe[28* 16 +: 16] = inputRe[14* 16 +: 16];
	assign fftIm[28* 16 +: 16] = inputIm[14* 16 +: 16];
	assign fftRe[29* 16 +: 16] = inputRe[46* 16 +: 16];
	assign fftIm[29* 16 +: 16] = inputIm[46* 16 +: 16];
	assign fftRe[30* 16 +: 16] = inputRe[30* 16 +: 16];
	assign fftIm[30* 16 +: 16] = inputIm[30* 16 +: 16];
	assign fftRe[31* 16 +: 16] = inputRe[62* 16 +: 16];
	assign fftIm[31* 16 +: 16] = inputIm[62* 16 +: 16];
	assign fftRe[32* 16 +: 16] = inputRe[1* 16 +: 16];
	assign fftIm[32* 16 +: 16] = inputIm[1* 16 +: 16];
	assign fftRe[33* 16 +: 16] = inputRe[33* 16 +: 16];
	assign fftIm[33* 16 +: 16] = inputIm[33* 16 +: 16];
	assign fftRe[34* 16 +: 16] = inputRe[17* 16 +: 16];
	assign fftIm[34* 16 +: 16] = inputIm[17* 16 +: 16];
	assign fftRe[35* 16 +: 16] = inputRe[49* 16 +: 16];
	assign fftIm[35* 16 +: 16] = inputIm[49* 16 +: 16];
	assign fftRe[36* 16 +: 16] = inputRe[9* 16 +: 16];
	assign fftIm[36* 16 +: 16] = inputIm[9* 16 +: 16];
	assign fftRe[37* 16 +: 16] = inputRe[41* 16 +: 16];
	assign fftIm[37* 16 +: 16] = inputIm[41* 16 +: 16];
	assign fftRe[38* 16 +: 16] = inputRe[25* 16 +: 16];
	assign fftIm[38* 16 +: 16] = inputIm[25* 16 +: 16];
	assign fftRe[39* 16 +: 16] = inputRe[57* 16 +: 16];
	assign fftIm[39* 16 +: 16] = inputIm[57* 16 +: 16];
	assign fftRe[40* 16 +: 16] = inputRe[5* 16 +: 16];
	assign fftIm[40* 16 +: 16] = inputIm[5* 16 +: 16];
	assign fftRe[41* 16 +: 16] = inputRe[37* 16 +: 16];
	assign fftIm[41* 16 +: 16] = inputIm[37* 16 +: 16];
	assign fftRe[42* 16 +: 16] = inputRe[21* 16 +: 16];
	assign fftIm[42* 16 +: 16] = inputIm[21* 16 +: 16];
	assign fftRe[43* 16 +: 16] = inputRe[53* 16 +: 16];
	assign fftIm[43* 16 +: 16] = inputIm[53* 16 +: 16];
	assign fftRe[44* 16 +: 16] = inputRe[13* 16 +: 16];
	assign fftIm[44* 16 +: 16] = inputIm[13* 16 +: 16];
	assign fftRe[45* 16 +: 16] = inputRe[45* 16 +: 16];
	assign fftIm[45* 16 +: 16] = inputIm[45* 16 +: 16];
	assign fftRe[46* 16 +: 16] = inputRe[29* 16 +: 16];
	assign fftIm[46* 16 +: 16] = inputIm[29* 16 +: 16];
	assign fftRe[47* 16 +: 16] = inputRe[61* 16 +: 16];
	assign fftIm[47* 16 +: 16] = inputIm[61* 16 +: 16];
	assign fftRe[48* 16 +: 16] = inputRe[3* 16 +: 15];
	assign fftIm[48* 16 +: 16] = inputIm[3* 16 +: 15];
	assign fftRe[49* 16 +: 16] = inputRe[35* 16 +: 16];
	assign fftIm[49* 16 +: 16] = inputIm[35* 16 +: 16];
	assign fftRe[50* 16 +: 16] = inputRe[19* 16 +: 16];
	assign fftIm[50* 16 +: 16] = inputIm[19* 16 +: 16];
	assign fftRe[51* 16 +: 16] = inputRe[51* 16 +: 16];
	assign fftIm[51* 16 +: 16] = inputIm[51* 16 +: 16];
	assign fftRe[52* 16 +: 16] = inputRe[11* 16 +: 16];
	assign fftIm[52* 16 +: 16] = inputIm[11* 16 +: 16];
	assign fftRe[53* 16 +: 16] = inputRe[43* 16 +: 16];
	assign fftIm[53* 16 +: 16] = inputIm[43* 16 +: 16];
	assign fftRe[54* 16 +: 16] = inputRe[27* 16 +: 16];
	assign fftIm[54* 16 +: 16] = inputIm[27* 16 +: 16];
	assign fftRe[55* 16 +: 16] = inputRe[59* 16 +: 16];
	assign fftIm[55* 16 +: 16] = inputIm[59* 16 +: 16];
	assign fftRe[56* 16 +: 16] = inputRe[7* 16 +: 15];
	assign fftIm[56* 16 +: 16] = inputIm[7* 16 +: 15];
	assign fftRe[57* 16 +: 16] = inputRe[39* 16 +: 16];
	assign fftIm[57* 16 +: 16] = inputIm[39* 16 +: 16];
	assign fftRe[58* 16 +: 16] = inputRe[23* 16 +: 16];
	assign fftIm[58* 16 +: 16] = inputIm[23* 16 +: 16];
	assign fftRe[59* 16 +: 16] = inputRe[55* 16 +: 16];
	assign fftIm[59* 16 +: 16] = inputIm[55* 16 +: 16];
	assign fftRe[60* 16 +: 16] = inputRe[15* 16 +: 16];
	assign fftIm[60* 16 +: 16] = inputIm[15* 16 +: 16];
	assign fftRe[61* 16 +: 16] = inputRe[47* 16 +: 16];
	assign fftIm[61* 16 +: 16] = inputIm[47* 16 +: 16];
	assign fftRe[62* 16 +: 16] = inputRe[31* 16 +: 16];
	assign fftIm[62* 16 +: 16] = inputIm[31* 16 +: 16];
	assign fftRe[63* 16 +: 16] = inputRe[63* 16 +: 16];
	assign fftIm[63* 16 +: 16] = inputIm[63* 16 +: 16];
	assign outputRe = fftRe;
	assign outputIm = fftIm;
endmodule
