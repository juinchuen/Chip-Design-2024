module InputSignalRouter #(
    parameter D_WIDTH = 64,
    parameter LOG_2_WIDTH = 6
) (
    input logic [15:0] inputRe [((D_WIDTH) - 1):0],
    input logic [15:0] inputIm [((D_WIDTH) - 1):0],
    output logic [15:0] outputRe [((D_WIDTH) - 1):0],
    output logic [15:0] outputIm [((D_WIDTH) - 1):0]
);
    // Correctly route the input signal

    logic [15:0] fftRe [((D_WIDTH) - 1):0];
    logic [15:0] fftIm [((D_WIDTH) - 1):0];
	assign fftRe[0] = inputRe[0];
	assign fftIm[0] = inputIm[0];
	assign fftRe[1] = inputRe[32];
	assign fftIm[1] = inputIm[32];
	assign fftRe[2] = inputRe[16];
	assign fftIm[2] = inputIm[16];
	assign fftRe[3] = inputRe[48];
	assign fftIm[3] = inputIm[48];
	assign fftRe[4] = inputRe[8];
	assign fftIm[4] = inputIm[8];
	assign fftRe[5] = inputRe[40];
	assign fftIm[5] = inputIm[40];
	assign fftRe[6] = inputRe[24];
	assign fftIm[6] = inputIm[24];
	assign fftRe[7] = inputRe[56];
	assign fftIm[7] = inputIm[56];
	assign fftRe[8] = inputRe[4];
	assign fftIm[8] = inputIm[4];
	assign fftRe[9] = inputRe[36];
	assign fftIm[9] = inputIm[36];
	assign fftRe[10] = inputRe[20];
	assign fftIm[10] = inputIm[20];
	assign fftRe[11] = inputRe[52];
	assign fftIm[11] = inputIm[52];
	assign fftRe[12] = inputRe[12];
	assign fftIm[12] = inputIm[12];
	assign fftRe[13] = inputRe[44];
	assign fftIm[13] = inputIm[44];
	assign fftRe[14] = inputRe[28];
	assign fftIm[14] = inputIm[28];
	assign fftRe[15] = inputRe[60];
	assign fftIm[15] = inputIm[60];
	assign fftRe[16] = inputRe[2];
	assign fftIm[16] = inputIm[2];
	assign fftRe[17] = inputRe[34];
	assign fftIm[17] = inputIm[34];
	assign fftRe[18] = inputRe[18];
	assign fftIm[18] = inputIm[18];
	assign fftRe[19] = inputRe[50];
	assign fftIm[19] = inputIm[50];
	assign fftRe[20] = inputRe[10];
	assign fftIm[20] = inputIm[10];
	assign fftRe[21] = inputRe[42];
	assign fftIm[21] = inputIm[42];
	assign fftRe[22] = inputRe[26];
	assign fftIm[22] = inputIm[26];
	assign fftRe[23] = inputRe[58];
	assign fftIm[23] = inputIm[58];
	assign fftRe[24] = inputRe[6];
	assign fftIm[24] = inputIm[6];
	assign fftRe[25] = inputRe[38];
	assign fftIm[25] = inputIm[38];
	assign fftRe[26] = inputRe[22];
	assign fftIm[26] = inputIm[22];
	assign fftRe[27] = inputRe[54];
	assign fftIm[27] = inputIm[54];
	assign fftRe[28] = inputRe[14];
	assign fftIm[28] = inputIm[14];
	assign fftRe[29] = inputRe[46];
	assign fftIm[29] = inputIm[46];
	assign fftRe[30] = inputRe[30];
	assign fftIm[30] = inputIm[30];
	assign fftRe[31] = inputRe[62];
	assign fftIm[31] = inputIm[62];
	assign fftRe[32] = inputRe[1];
	assign fftIm[32] = inputIm[1];
	assign fftRe[33] = inputRe[33];
	assign fftIm[33] = inputIm[33];
	assign fftRe[34] = inputRe[17];
	assign fftIm[34] = inputIm[17];
	assign fftRe[35] = inputRe[49];
	assign fftIm[35] = inputIm[49];
	assign fftRe[36] = inputRe[9];
	assign fftIm[36] = inputIm[9];
	assign fftRe[37] = inputRe[41];
	assign fftIm[37] = inputIm[41];
	assign fftRe[38] = inputRe[25];
	assign fftIm[38] = inputIm[25];
	assign fftRe[39] = inputRe[57];
	assign fftIm[39] = inputIm[57];
	assign fftRe[40] = inputRe[5];
	assign fftIm[40] = inputIm[5];
	assign fftRe[41] = inputRe[37];
	assign fftIm[41] = inputIm[37];
	assign fftRe[42] = inputRe[21];
	assign fftIm[42] = inputIm[21];
	assign fftRe[43] = inputRe[53];
	assign fftIm[43] = inputIm[53];
	assign fftRe[44] = inputRe[13];
	assign fftIm[44] = inputIm[13];
	assign fftRe[45] = inputRe[45];
	assign fftIm[45] = inputIm[45];
	assign fftRe[46] = inputRe[29];
	assign fftIm[46] = inputIm[29];
	assign fftRe[47] = inputRe[61];
	assign fftIm[47] = inputIm[61];
	assign fftRe[48] = inputRe[3];
	assign fftIm[48] = inputIm[3];
	assign fftRe[49] = inputRe[35];
	assign fftIm[49] = inputIm[35];
	assign fftRe[50] = inputRe[19];
	assign fftIm[50] = inputIm[19];
	assign fftRe[51] = inputRe[51];
	assign fftIm[51] = inputIm[51];
	assign fftRe[52] = inputRe[11];
	assign fftIm[52] = inputIm[11];
	assign fftRe[53] = inputRe[43];
	assign fftIm[53] = inputIm[43];
	assign fftRe[54] = inputRe[27];
	assign fftIm[54] = inputIm[27];
	assign fftRe[55] = inputRe[59];
	assign fftIm[55] = inputIm[59];
	assign fftRe[56] = inputRe[7];
	assign fftIm[56] = inputIm[7];
	assign fftRe[57] = inputRe[39];
	assign fftIm[57] = inputIm[39];
	assign fftRe[58] = inputRe[23];
	assign fftIm[58] = inputIm[23];
	assign fftRe[59] = inputRe[55];
	assign fftIm[59] = inputIm[55];
	assign fftRe[60] = inputRe[15];
	assign fftIm[60] = inputIm[15];
	assign fftRe[61] = inputRe[47];
	assign fftIm[61] = inputIm[47];
	assign fftRe[62] = inputRe[31];
	assign fftIm[62] = inputIm[31];
	assign fftRe[63] = inputRe[63];
	assign fftIm[63] = inputIm[63];
	assign outputRe = fftRe;
	assign outputIm = fftIm;
endmodule
